//instance를 배우는 코드임

module top_module ( input a, input b, output out );
    mod_a instance_name (.out(out), .in1(a), .in2(b));
endmodule